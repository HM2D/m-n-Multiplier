module or65(out,a,b);
input [64:0] a,b;
output [64:0] out;

assign out = a|b;

endmodule
