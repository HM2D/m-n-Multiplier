module not65(out,a);
input [64:0] a;
output wire [64:0] out;

assign out = ~a;

endmodule


